`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:58:48 02/25/2015 
// Design Name: 
// Module Name:    IM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module IM(
    input [7:0] Address,
    output wire [31:0] InstructionOut
    );
	 
	 reg [31:0] iM [255:0];
	 
	 assign InstructionOut = iM[Address[7:0]];
	 
	 initial begin
		
		//iM[0] = 8'h8c;
		//iM[1] = 8'h05;
		//iM[2] = 8'h14;
		//iM[3] = 8'h8c;
		//iM[4] = 8'h0a;
		//iM[5] = 8'h14;
	


	
		iM[0] = 32'b 100011_00000_00101_0000000000010100;
		iM[1] = 32'b 100011_00000_00101_0000000000010100;
		iM[2] = 32'b 100011_00000_00101_0000000000010100;
		iM[3] = 32'b 100011_00000_00101_0000000000010100;
		iM[4] = 32'b 100011_00000_00101_0000000000010100;
		iM[5] = 32'b 100011_00000_00101_0000000000010100;
		iM[6] = 32'b 100011_00000_00101_0000000000010100;
		iM[7] = 32'b 100011_00000_00101_0000000000010100;

		iM[20] = 32'b 100011_00000_00101_0000000000010100; 
		iM[21] = 32'b 100011_00000_00101_0000000000010100;
		iM[22] = 32'b 100011_00000_00101_0000000000010100;
		iM[23] = 32'b 100011_00000_00101_0000000000010100;

		iM[40] = 32'b 100011_00000_00101_0000000000010100;
		iM[41] = 32'b 100011_00000_00101_0000000000010100;
		iM[42] = 32'b 100011_00000_00101_0000000000010100;
		iM[43] = 32'b 100011_00000_00101_0000000000010100;

	end	 
	 


endmodule
